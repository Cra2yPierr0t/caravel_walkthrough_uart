rggen-verilog-rtl/rggen_rtl_macros.vh